class AES_TEST;
    
    
    
endclass
