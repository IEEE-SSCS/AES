class fill;
bit[127:0] katvk[bit[127:0]];
bit[127:0] katvt [bit[127:0]];
  task  fill; 
    
   katvt='{
128'h80000000000000000000000000000000	: 128'h3ad78e726c1ec02b7ebfe92b23d9ec34,
128'hc0000000000000000000000000000000	: 128'haae5939c8efdf2f04e60b9fe7117b2c2,
128'he0000000000000000000000000000000	: 128'hf031d4d74f5dcbf39daaf8ca3af6e527,
128'hf0000000000000000000000000000000	: 128'h96d9fd5cc4f07441727df0f33e401a36,
128'hf8000000000000000000000000000000	: 128'h30ccdb044646d7e1f3ccea3dca08b8c0,
128'hfc000000000000000000000000000000	: 128'h16ae4ce5042a67ee8e177b7c587ecc82,
128'hfe000000000000000000000000000000	: 128'hb6da0bb11a23855d9c5cb1b4c6412e0a,
128'hff000000000000000000000000000000	: 128'hdb4f1aa530967d6732ce4715eb0ee24b,
128'hff800000000000000000000000000000	: 128'ha81738252621dd180a34f3455b4baa2f,
128'hffc00000000000000000000000000000	: 128'h77e2b508db7fd89234caf7939ee5621a,
128'hffe00000000000000000000000000000	: 128'hb8499c251f8442ee13f0933b688fcd19,
128'hfff00000000000000000000000000000	: 128'h965135f8a81f25c9d630b17502f68e53,
128'hfff80000000000000000000000000000	: 128'h8b87145a01ad1c6cede995ea3670454f,
128'hfffc0000000000000000000000000000	: 128'h8eae3b10a0c8ca6d1d3b0fa61e56b0b2,
128'hfffc0000000000000000000000000000	: 128'h8eae3b10a0c8ca6d1d3b0fa61e56b0b2,
128'hfffe0000000000000000000000000000	: 128'h64b4d629810fda6bafdf08f3b0d8d2c5,
128'hffff0000000000000000000000000000	: 128'hd7e5dbd3324595f8fdc7d7c571da6c2a,
128'hffff8000000000000000000000000000	: 128'hf3f72375264e167fca9de2c1527d9606,
128'hffffc000000000000000000000000000	: 128'h8ee79dd4f401ff9b7ea945d86666c13b,
128'hffffe000000000000000000000000000	: 128'hdd35cea2799940b40db3f819cb94c08b,
128'hfffff000000000000000000000000000	: 128'h6941cb6b3e08c2b7afa581ebdd607b87,
128'hfffff800000000000000000000000000	: 128'h2c20f439f6bb097b29b8bd6d99aad799,
128'hfffffc00000000000000000000000000	: 128'h625d01f058e565f77ae86378bd2c49b3,
128'hfffffe00000000000000000000000000	: 128'hc0b5fd98190ef45fbb4301438d095950,
128'hffffff00000000000000000000000000	: 128'h13001ff5d99806efd25da34f56be854b,
128'hffffff80000000000000000000000000	: 128'h3b594c60f5c8277a5113677f94208d82,
128'hffffffc0000000000000000000000000	: 128'he9c0fc1818e4aa46bd2e39d638f89e05,
128'hffffffe0000000000000000000000000	: 128'hf8023ee9c3fdc45a019b4e985c7e1a54,
128'hfffffff0000000000000000000000000	: 128'h35f40182ab4662f3023baec1ee796b57,
128'hfffffff8000000000000000000000000	: 128'h3aebbad7303649b4194a6945c6cc3694,
128'hfffffffc000000000000000000000000	: 128'ha2124bea53ec2834279bed7f7eb0f938,
128'hfffffffe000000000000000000000000	: 128'hb9fb4399fa4facc7309e14ec98360b0a,
128'hffffffff000000000000000000000000	: 128'hc26277437420c5d634f715aea81a9132,
128'hffffffff800000000000000000000000	: 128'h171a0e1b2dd424f0e089af2c4c10f32f,
128'hffffffffc00000000000000000000000	: 128'h7cadbe402d1b208fe735edce00aee7ce,
128'hffffffffe00000000000000000000000	: 128'h43b02ff929a1485af6f5c6d6558baa0f,
128'hfffffffff00000000000000000000000	: 128'h092faacc9bf43508bf8fa8613ca75dea,
128'hfffffffff80000000000000000000000	: 128'hcb2bf8280f3f9742c7ed513fe802629c,
128'hfffffffffc0000000000000000000000	: 128'h215a41ee442fa992a6e323986ded3f68,
128'hfffffffffe0000000000000000000000	: 128'hf21e99cf4f0f77cea836e11a2fe75fb1,
128'hffffffffff0000000000000000000000	: 128'h95e3a0ca9079e646331df8b4e70d2cd6,
128'hffffffffff8000000000000000000000	: 128'h4afe7f120ce7613f74fc12a01a828073,
128'hffffffffffc000000000000000000000	: 128'h827f000e75e2c8b9d479beed913fe678,
128'hffffffffffe000000000000000000000	: 128'h35830c8e7aaefe2d30310ef381cbf691,
128'hfffffffffff000000000000000000000	: 128'h191aa0f2c8570144f38657ea4085ebe5,
128'hfffffffffff800000000000000000000	: 128'h85062c2c909f15d9269b6c18ce99c4f0,
128'hfffffffffffc00000000000000000000	: 128'h678034dc9e41b5a560ed239eeab1bc78,
128'hfffffffffffe00000000000000000000	: 128'hc2f93a4ce5ab6d5d56f1b93cf19911c1,
128'hffffffffffff00000000000000000000	: 128'h1c3112bcb0c1dcc749d799743691bf82,
128'hffffffffffff80000000000000000000	: 128'h00c55bd75c7f9c881989d3ec1911c0d4,
128'hffffffffffffc0000000000000000000	: 128'hea2e6b5ef182b7dff3629abd6a12045f,
128'hffffffffffffe0000000000000000000	: 128'h22322327e01780b17397f24087f8cc6f,
128'hfffffffffffff0000000000000000000	: 128'hc9cacb5cd11692c373b2411768149ee7,
128'hfffffffffffff8000000000000000000	: 128'ha18e3dbbca577860dab6b80da3139256,
128'hfffffffffffffc000000000000000000	: 128'h79b61c37bf328ecca8d743265a3d425c,
128'hfffffffffffffe000000000000000000	: 128'hd2d99c6bcc1f06fda8e27e8ae3f1ccc7,
128'hffffffffffffff000000000000000000	: 128'h1bfd4b91c701fd6b61b7f997829d663b,
128'hffffffffffffff800000000000000000	: 128'h11005d52f25f16bdc9545a876a63490a,
128'hffffffffffffffc00000000000000000	: 128'h3a4d354f02bb5a5e47d39666867f246a,
128'hffffffffffffffe00000000000000000	: 128'hd451b8d6e1e1a0ebb155fbbf6e7b7dc3,
128'hfffffffffffffff00000000000000000	: 128'h6898d4f42fa7ba6a10ac05e87b9f2080,
128'hfffffffffffffff80000000000000000	: 128'hb611295e739ca7d9b50f8e4c0e754a3f,
128'hfffffffffffffffc0000000000000000	: 128'h7d33fc7d8abe3ca1936759f8f5deaf20,
128'hfffffffffffffffe0000000000000000	: 128'h3b5e0f566dc96c298f0c12637539b25c,
128'hffffffffffffffff0000000000000000	: 128'hf807c3e7985fe0f5a50e2cdb25c5109e,
128'hffffffffffffffff8000000000000000	: 128'h41f992a856fb278b389a62f5d274d7e9,
128'hffffffffffffffffc000000000000000	: 128'h10d3ed7a6fe15ab4d91acbc7d0767ab1,
128'hffffffffffffffffe000000000000000	: 128'h21feecd45b2e675973ac33bf0c5424fc,
128'hfffffffffffffffff000000000000000	: 128'h1480cb3955ba62d09eea668f7c708817,
128'hfffffffffffffffff800000000000000	: 128'h66404033d6b72b609354d5496e7eb511,
128'hfffffffffffffffffc00000000000000	: 128'h1c317a220a7d700da2b1e075b00266e1,
128'hfffffffffffffffffe00000000000000	: 128'hab3b89542233f1271bf8fd0c0f403545,
128'hffffffffffffffffff00000000000000	: 128'hd93eae966fac46dca927d6b114fa3f9e,
128'hffffffffffffffffff80000000000000	: 128'h1bdec521316503d9d5ee65df3ea94ddf,
128'hffffffffffffffffffc0000000000000	: 128'heef456431dea8b4acf83bdae3717f75f,
128'hffffffffffffffffffe0000000000000	: 128'h06f2519a2fafaa596bfef5cfa15c21b9,
128'hfffffffffffffffffff0000000000000	: 128'h251a7eac7e2fe809e4aa8d0d7012531a,
128'hfffffffffffffffffff8000000000000	: 128'h3bffc16e4c49b268a20f8d96a60b4058,
128'hfffffffffffffffffffc000000000000	: 128'he886f9281999c5bb3b3e8862e2f7c988,
128'hfffffffffffffffffffe000000000000	: 128'h563bf90d61beef39f48dd625fcef1361,
128'hffffffffffffffffffff000000000000	: 128'h4d37c850644563c69fd0acd9a049325b,
128'hffffffffffffffffffff800000000000	: 128'hb87c921b91829ef3b13ca541ee1130a6,
128'hffffffffffffffffffffc00000000000	: 128'h2e65eb6b6ea383e109accce8326b0393,
128'hffffffffffffffffffffe00000000000	: 128'h9ca547f7439edc3e255c0f4d49aa8990,
128'hfffffffffffffffffffff00000000000	: 128'ha5e652614c9300f37816b1f9fd0c87f9,
128'hfffffffffffffffffffff80000000000	: 128'h14954f0b4697776f44494fe458d814ed,
128'hfffffffffffffffffffffc0000000000	: 128'h7c8d9ab6c2761723fe42f8bb506cbcf7,
128'hfffffffffffffffffffffe0000000000	: 128'hdb7e1932679fdd99742aab04aa0d5a80,
128'hffffffffffffffffffffff0000000000	: 128'h4c6a1c83e568cd10f27c2d73ded19c28,
128'hffffffffffffffffffffff8000000000	: 128'h90ecbe6177e674c98de412413f7ac915,
128'hffffffffffffffffffffffc000000000	: 128'h90684a2ac55fe1ec2b8ebd5622520b73,
128'hffffffffffffffffffffffe000000000	: 128'h7472f9a7988607ca79707795991035e6,
128'hfffffffffffffffffffffff000000000	: 128'h56aff089878bf3352f8df172a3ae47d8,
128'hfffffffffffffffffffffff800000000	: 128'h65c0526cbe40161b8019a2a3171abd23,
128'hfffffffffffffffffffffffc00000000	: 128'h377be0be33b4e3e310b4aabda173f84f,
128'hfffffffffffffffffffffffe00000000	: 128'h9402e9aa6f69de6504da8d20c4fcaa2f,
128'hffffffffffffffffffffffff00000000	: 128'h123c1f4af313ad8c2ce648b2e71fb6e1,
128'hffffffffffffffffffffffff80000000	: 128'h1ffc626d30203dcdb0019fb80f726cf4,
128'hffffffffffffffffffffffffc0000000	: 128'h76da1fbe3a50728c50fd2e621b5ad885,
128'hffffffffffffffffffffffffe0000000	: 128'h082eb8be35f442fb52668e16a591d1d6,
128'hfffffffffffffffffffffffff0000000	: 128'he656f9ecf5fe27ec3e4a73d00c282fb3,
128'hfffffffffffffffffffffffff8000000	: 128'h2ca8209d63274cd9a29bb74bcd77683a,
128'hfffffffffffffffffffffffffc000000	: 128'h79bf5dce14bb7dd73a8e3611de7ce026,
128'hfffffffffffffffffffffffffe000000	: 128'h3c849939a5d29399f344c4a0eca8a576,
128'hffffffffffffffffffffffffff000000	: 128'hed3c0a94d59bece98835da7aa4f07ca2,
128'hffffffffffffffffffffffffff800000	: 128'h63919ed4ce10196438b6ad09d99cd795,
128'hffffffffffffffffffffffffffc00000	: 128'h7678f3a833f19fea95f3c6029e2bc610,
128'hffffffffffffffffffffffffffe00000	: 128'h3aa426831067d36b92be7c5f81c13c56,
128'hfffffffffffffffffffffffffff00000	: 128'h9272e2d2cdd11050998c845077a30ea0,
128'hfffffffffffffffffffffffffff80000	: 128'h088c4b53f5ec0ff814c19adae7f6246c,
128'hfffffffffffffffffffffffffffc0000	: 128'h4010a5e401fdf0a0354ddbcc0d012b17,
128'hfffffffffffffffffffffffffffe0000	: 128'ha87a385736c0a6189bd6589bd8445a93,
128'hffffffffffffffffffffffffffff0000	: 128'h545f2b83d9616dccf60fa9830e9cd287,
128'hffffffffffffffffffffffffffff8000	: 128'h4b706f7f92406352394037a6d4f4688d,
128'hffffffffffffffffffffffffffffc000	: 128'hb7972b3941c44b90afa7b264bfba7387,
128'hffffffffffffffffffffffffffffe000	: 128'h6f45732cf10881546f0fd23896d2bb60,
128'hfffffffffffffffffffffffffffff000	: 128'h2e3579ca15af27f64b3c955a5bfc30ba,
128'hfffffffffffffffffffffffffffff800	: 128'h34a2c5a91ae2aec99b7d1b5fa6780447,
128'hfffffffffffffffffffffffffffffc00	: 128'ha4d6616bd04f87335b0e53351227a9ee,
128'hfffffffffffffffffffffffffffffe00	: 128'h7f692b03945867d16179a8cefc83ea3f,
128'hffffffffffffffffffffffffffffff00	: 128'h3bd141ee84a0e6414a26e7a4f281f8a2,
128'hffffffffffffffffffffffffffffff80	: 128'hd1788f572d98b2b16ec5d5f3922b99bc,
128'hffffffffffffffffffffffffffffffc0	: 128'h0833ff6f61d98a57b288e8c3586b85a6,
128'hffffffffffffffffffffffffffffffe0	: 128'h8568261797de176bf0b43becc6285afb,
128'hfffffffffffffffffffffffffffffff0	: 128'hf9b0fda0c4a898f5b9e6f661c4ce4d07,
128'hfffffffffffffffffffffffffffffff8	: 128'h8ade895913685c67c5269f8aae42983e,
128'hfffffffffffffffffffffffffffffffc	: 128'h39bde67d5c8ed8a8b1c37eb8fa9f5ac0,
128'hfffffffffffffffffffffffffffffffe	: 128'h5c005e72c1418c44f569f2ea33ba54f3,
128'hffffffffffffffffffffffffffffffff	: 128'h3f5b8cc9ea855a0afa7347d23e8d664e
};
   katvk='{
128'h80000000000000000000000000000000	: 128'h0edd33d3c621e546455bd8ba1418bec8,
128'hc0000000000000000000000000000000	: 128'h4bc3f883450c113c64ca42e1112a9e87,
128'he0000000000000000000000000000000	: 128'h72a1da770f5d7ac4c9ef94d822affd97,
128'hf0000000000000000000000000000000	: 128'h970014d634e2b7650777e8e84d03ccd8,
128'hf8000000000000000000000000000000	: 128'hf17e79aed0db7e279e955b5f493875a7,
128'hfc000000000000000000000000000000	: 128'h9ed5a75136a940d0963da379db4af26a,
128'hfe000000000000000000000000000000	: 128'hc4295f83465c7755e8fa364bac6a7ea5,
128'hff000000000000000000000000000000	: 128'hb1d758256b28fd850ad4944208cf1155,
128'hff800000000000000000000000000000	: 128'h42ffb34c743de4d88ca38011c990890b,
128'hffc00000000000000000000000000000	: 128'h9958f0ecea8b2172c0c1995f9182c0f3,
128'hffe00000000000000000000000000000	: 128'h956d7798fac20f82a8823f984d06f7f5,
128'hfff00000000000000000000000000000	: 128'ha01bf44f2d16be928ca44aaf7b9b106b,
128'hfff80000000000000000000000000000	: 128'hb5f1a33e50d40d103764c76bd4c6b6f8,
128'hfffc0000000000000000000000000000	: 128'h2637050c9fc0d4817e2d69de878aee8d,
128'hfffe0000000000000000000000000000	: 128'h113ecbe4a453269a0dd26069467fb5b5,
128'hffff0000000000000000000000000000	: 128'h97d0754fe68f11b9e375d070a608c884,
128'hffff8000000000000000000000000000	: 128'hc6a0b3e998d05068a5399778405200b4,
128'hffffc000000000000000000000000000	: 128'hdf556a33438db87bc41b1752c55e5e49,
128'hffffe000000000000000000000000000	: 128'h90fb128d3a1af6e548521bb962bf1f05,
128'hfffff000000000000000000000000000	: 128'h26298e9c1db517c215fadfb7d2a8d691,
128'hfffff800000000000000000000000000	: 128'ha6cb761d61f8292d0df393a279ad0380,
128'hfffffc00000000000000000000000000	: 128'h12acd89b13cd5f8726e34d44fd486108,
128'hfffffe00000000000000000000000000	: 128'h95b1703fc57ba09fe0c3580febdd7ed4,
128'hffffff00000000000000000000000000	: 128'hde11722d893e9f9121c381becc1da59a,
128'hffffff80000000000000000000000000	: 128'h6d114ccb27bf391012e8974c546d9bf2,
128'hffffffc0000000000000000000000000	: 128'h5ce37e17eb4646ecfac29b9cc38d9340,
128'hffffffe0000000000000000000000000	: 128'h18c1b6e2157122056d0243d8a165cddb,
128'hfffffff0000000000000000000000000	: 128'h99693e6a59d1366c74d823562d7e1431,
128'hfffffff8000000000000000000000000	: 128'h6c7c64dc84a8bba758ed17eb025a57e3,
128'hfffffffc000000000000000000000000	: 128'he17bc79f30eaab2fac2cbbe3458d687a,
128'hfffffffe000000000000000000000000	: 128'h1114bc2028009b923f0b01915ce5e7c4,
128'hffffffff000000000000000000000000	: 128'h9c28524a16a1e1c1452971caa8d13476,
128'hffffffff800000000000000000000000	: 128'hed62e16363638360fdd6ad62112794f0,
128'hffffffffc00000000000000000000000	: 128'h5a8688f0b2a2c16224c161658ffd4044,
128'hffffffffe00000000000000000000000	: 128'h23f710842b9bb9c32f26648c786807ca,
128'hfffffffff00000000000000000000000	: 128'h44a98bf11e163f632c47ec6a49683a89,
128'hfffffffff80000000000000000000000	: 128'h0f18aff94274696d9b61848bd50ac5e5,
128'hfffffffffc0000000000000000000000	: 128'h82408571c3e2424540207f833b6dda69,
128'hfffffffffe0000000000000000000000	: 128'h303ff996947f0c7d1f43c8f3027b9b75,
128'hffffffffff0000000000000000000000	: 128'h7df4daf4ad29a3615a9b6ece5c99518a,
128'hffffffffff8000000000000000000000	: 128'hc72954a48d0774db0b4971c526260415,
128'hffffffffffc000000000000000000000	: 128'h1df9b76112dc6531e07d2cfda04411f0,
128'hffffffffffe000000000000000000000	: 128'h8e4d8e699119e1fc87545a647fb1d34f,
128'hfffffffffff000000000000000000000	: 128'he6c4807ae11f36f091c57d9fb68548d1,
128'hfffffffffff800000000000000000000	: 128'h8ebf73aad49c82007f77a5c1ccec6ab4,
128'hfffffffffffc00000000000000000000	: 128'h4fb288cc2040049001d2c7585ad123fc,
128'hfffffffffffe00000000000000000000	: 128'h04497110efb9dceb13e2b13fb4465564,
128'hffffffffffff00000000000000000000	: 128'h75550e6cb5a88e49634c9ab69eda0430,
128'hffffffffffff80000000000000000000	: 128'hb6768473ce9843ea66a81405dd50b345,
128'hffffffffffffc0000000000000000000	: 128'hcb2f430383f9084e03a653571e065de6,
128'hffffffffffffe0000000000000000000	: 128'hff4e66c07bae3e79fb7d210847a3b0ba,
128'hfffffffffffff0000000000000000000	: 128'h7b90785125505fad59b13c186dd66ce3,
128'hfffffffffffff8000000000000000000	: 128'h8b527a6aebdaec9eaef8eda2cb7783e5,
128'hfffffffffffffc000000000000000000	: 128'h43fdaf53ebbc9880c228617d6a9b548b,
128'hfffffffffffffe000000000000000000	: 128'h53786104b9744b98f052c46f1c850d0b,
128'hffffffffffffff000000000000000000	: 128'hb5ab3013dd1e61df06cbaf34ca2aee78,
128'hffffffffffffff800000000000000000	: 128'h7470469be9723030fdcc73a8cd4fbb10,
128'hffffffffffffffc00000000000000000	: 128'ha35a63f5343ebe9ef8167bcb48ad122e,
128'hffffffffffffffe00000000000000000	: 128'hfd8687f0757a210e9fdf181204c30863,
128'hfffffffffffffff00000000000000000	: 128'h7a181e84bd5457d26a88fbae96018fb0,
128'hfffffffffffffff80000000000000000	: 128'h653317b9362b6f9b9e1a580e68d494b5,
128'hfffffffffffffffc0000000000000000	: 128'h995c9dc0b689f03c45867b5faa5c18d1,
128'hfffffffffffffffe0000000000000000	: 128'h77a4d96d56dda398b9aabecfc75729fd,
128'hffffffffffffffff0000000000000000	: 128'h84be19e053635f09f2665e7bae85b42d,
128'hffffffffffffffff8000000000000000	: 128'h32cd652842926aea4aa6137bb2be2b5e,
128'hffffffffffffffffc000000000000000	: 128'h493d4a4f38ebb337d10aa84e9171a554,
128'hffffffffffffffffe000000000000000	: 128'hd9bff7ff454b0ec5a4a2a69566e2cb84,
128'hfffffffffffffffff000000000000000	: 128'h3535d565ace3f31eb249ba2cc6765d7a,
128'hfffffffffffffffff800000000000000	: 128'hf60e91fc3269eecf3231c6e9945697c6,
128'hfffffffffffffffffc00000000000000	: 128'hab69cfadf51f8e604d9cc37182f6635a,
128'hfffffffffffffffffe00000000000000	: 128'h7866373f24a0b6ed56e0d96fcdafb877,
128'hffffffffffffffffff00000000000000	: 128'h1ea448c2aac954f5d812e9d78494446a,
128'hffffffffffffffffff80000000000000	: 128'hacc5599dd8ac02239a0fef4a36dd1668,
128'hffffffffffffffffffc0000000000000	: 128'hd8764468bb103828cf7e1473ce895073,
128'hffffffffffffffffffe0000000000000	: 128'h1b0d02893683b9f180458e4aa6b73982,
128'hfffffffffffffffffff0000000000000	: 128'h96d9b017d302df410a937dcdb8bb6e43,
128'hfffffffffffffffffff8000000000000	: 128'hef1623cc44313cff440b1594a7e21cc6,
128'hfffffffffffffffffffc000000000000	: 128'h284ca2fa35807b8b0ae4d19e11d7dbd7,
128'hfffffffffffffffffffe000000000000	: 128'hf2e976875755f9401d54f36e2a23a594,
128'hffffffffffffffffffff000000000000	: 128'hec198a18e10e532403b7e20887c8dd80,
128'hffffffffffffffffffff800000000000	: 128'h545d50ebd919e4a6949d96ad47e46a80,
128'hffffffffffffffffffffc00000000000	: 128'hdbdfb527060e0a71009c7bb0c68f1d44,
128'hffffffffffffffffffffe00000000000	: 128'h9cfa1322ea33da2173a024f2ff0d896d,
128'hfffffffffffffffffffff00000000000	: 128'h8785b1a75b0f3bd958dcd0e29318c521,
128'hfffffffffffffffffffff80000000000	: 128'h38f67b9e98e4a97b6df030a9fcdd0104,
128'hfffffffffffffffffffffc0000000000	: 128'h192afffb2c880e82b05926d0fc6c448b,
128'hfffffffffffffffffffffe0000000000	: 128'h6a7980ce7b105cf530952d74daaf798c,
128'hffffffffffffffffffffff0000000000	: 128'hea3695e1351b9d6858bd958cf513ef6c,
128'hffffffffffffffffffffff8000000000	: 128'h6da0490ba0ba0343b935681d2cce5ba1,
128'hffffffffffffffffffffffc000000000	: 128'hf0ea23af08534011c60009ab29ada2f1,
128'hffffffffffffffffffffffe000000000	: 128'hff13806cf19cc38721554d7c0fcdcd4b,
128'hfffffffffffffffffffffff000000000	: 128'h6838af1f4f69bae9d85dd188dcdf0688,
128'hfffffffffffffffffffffff800000000	: 128'h36cf44c92d550bfb1ed28ef583ddf5d7,
128'hfffffffffffffffffffffffc00000000	: 128'hd06e3195b5376f109d5c4ec6c5d62ced,
128'hfffffffffffffffffffffffe00000000	: 128'hc440de014d3d610707279b13242a5c36,
128'hffffffffffffffffffffffff00000000	: 128'hf0c5c6ffa5e0bd3a94c88f6b6f7c16b9,
128'hffffffffffffffffffffffff80000000	: 128'h3e40c3901cd7effc22bffc35dee0b4d9,
128'hffffffffffffffffffffffffc0000000	: 128'hb63305c72bedfab97382c406d0c49bc6,
128'hffffffffffffffffffffffffe0000000	: 128'h36bbaab22a6bd4925a99a2b408d2dbae,
128'hfffffffffffffffffffffffff0000000	: 128'h307c5b8fcd0533ab98bc51e27a6ce461,
128'hfffffffffffffffffffffffff8000000	: 128'h829c04ff4c07513c0b3ef05c03e337b5,
128'hfffffffffffffffffffffffffc000000	: 128'hf17af0e895dda5eb98efc68066e84c54,
128'hfffffffffffffffffffffffffe000000	: 128'h277167f3812afff1ffacb4a934379fc3,
128'hffffffffffffffffffffffffff000000	: 128'h2cb1dc3a9c72972e425ae2ef3eb597cd,
128'hffffffffffffffffffffffffff800000	: 128'h36aeaa3a213e968d4b5b679d3a2c97fe,
128'hffffffffffffffffffffffffffc00000	: 128'h9241daca4fdd034a82372db50e1a0f3f,
128'hffffffffffffffffffffffffffe00000	: 128'hc14574d9cd00cf2b5a7f77e53cd57885,
128'hfffffffffffffffffffffffffff00000	: 128'h793de39236570aba83ab9b737cb521c9,
128'hfffffffffffffffffffffffffff80000	: 128'h16591c0f27d60e29b85a96c33861a7ef,
128'hfffffffffffffffffffffffffffc0000	: 128'h44fb5c4d4f5cb79be5c174a3b1c97348,
128'hfffffffffffffffffffffffffffe0000	: 128'h674d2b61633d162be59dde04222f4740,
128'hffffffffffffffffffffffffffff0000	: 128'hb4750ff263a65e1f9e924ccfd98f3e37,
128'hffffffffffffffffffffffffffff8000	: 128'h62d0662d6eaeddedebae7f7ea3a4f6b6,
128'hffffffffffffffffffffffffffffc000	: 128'h70c46bb30692be657f7eaa93ebad9897,
128'hffffffffffffffffffffffffffffe000	: 128'h323994cfb9da285a5d9642e1759b224a,
128'hfffffffffffffffffffffffffffff000	: 128'h1dbf57877b7b17385c85d0b54851e371,
128'hfffffffffffffffffffffffffffff800	: 128'hdfa5c097cdc1532ac071d57b1d28d1bd,
128'hfffffffffffffffffffffffffffffc00	: 128'h3a0c53fa37311fc10bd2a9981f513174,
128'hfffffffffffffffffffffffffffffe00	: 128'hba4f970c0a25c41814bdae2e506be3b4,
128'hffffffffffffffffffffffffffffff00	: 128'h2dce3acb727cd13ccd76d425ea56e4f6,
128'hffffffffffffffffffffffffffffff80	: 128'h5160474d504b9b3eefb68d35f245f4b3,
128'hffffffffffffffffffffffffffffffc0	: 128'h41a8a947766635dec37553d9a6c0cbb7,
128'hffffffffffffffffffffffffffffffe0	: 128'h25d6cfe6881f2bf497dd14cd4ddf445b,
128'hfffffffffffffffffffffffffffffff0	: 128'h41c78c135ed9e98c096640647265da1e,
128'hfffffffffffffffffffffffffffffff8	: 128'h5a4d404d8917e353e92a21072c3b2305,
128'hfffffffffffffffffffffffffffffffc	: 128'h02bc96846b3fdc71643f384cd3cc3eaf,
128'hfffffffffffffffffffffffffffffffe	: 128'h9ba4a9143f4e5d4048521c4f8877d88e,
128'hffffffffffffffffffffffffffffffff	: 128'ha1f6258c877d5fcd8964484538bfc92c
};
  endtask
endclass 