class AES_test;
      
    
    
    
endclass
